module registerFile(
  input         clock,
  input         reset,
  input         io_regWrite,
  input  [4:0]  io_rs1_sel,
  input  [4:0]  io_rs2_sel,
  input  [4:0]  io_rd_sel,
  input  [31:0] io_writeData,
  output [31:0] io_rs1,
  output [31:0] io_rs2
);
  reg [31:0] registers_0; // @[registerFile.scala 15:26]
  reg [31:0] _RAND_0;
  reg [31:0] registers_1; // @[registerFile.scala 15:26]
  reg [31:0] _RAND_1;
  reg [31:0] registers_2; // @[registerFile.scala 15:26]
  reg [31:0] _RAND_2;
  reg [31:0] registers_3; // @[registerFile.scala 15:26]
  reg [31:0] _RAND_3;
  reg [31:0] registers_4; // @[registerFile.scala 15:26]
  reg [31:0] _RAND_4;
  reg [31:0] registers_5; // @[registerFile.scala 15:26]
  reg [31:0] _RAND_5;
  reg [31:0] registers_6; // @[registerFile.scala 15:26]
  reg [31:0] _RAND_6;
  reg [31:0] registers_7; // @[registerFile.scala 15:26]
  reg [31:0] _RAND_7;
  reg [31:0] registers_8; // @[registerFile.scala 15:26]
  reg [31:0] _RAND_8;
  reg [31:0] registers_9; // @[registerFile.scala 15:26]
  reg [31:0] _RAND_9;
  reg [31:0] registers_10; // @[registerFile.scala 15:26]
  reg [31:0] _RAND_10;
  reg [31:0] registers_11; // @[registerFile.scala 15:26]
  reg [31:0] _RAND_11;
  reg [31:0] registers_12; // @[registerFile.scala 15:26]
  reg [31:0] _RAND_12;
  reg [31:0] registers_13; // @[registerFile.scala 15:26]
  reg [31:0] _RAND_13;
  reg [31:0] registers_14; // @[registerFile.scala 15:26]
  reg [31:0] _RAND_14;
  reg [31:0] registers_15; // @[registerFile.scala 15:26]
  reg [31:0] _RAND_15;
  reg [31:0] registers_16; // @[registerFile.scala 15:26]
  reg [31:0] _RAND_16;
  reg [31:0] registers_17; // @[registerFile.scala 15:26]
  reg [31:0] _RAND_17;
  reg [31:0] registers_18; // @[registerFile.scala 15:26]
  reg [31:0] _RAND_18;
  reg [31:0] registers_19; // @[registerFile.scala 15:26]
  reg [31:0] _RAND_19;
  reg [31:0] registers_20; // @[registerFile.scala 15:26]
  reg [31:0] _RAND_20;
  reg [31:0] registers_21; // @[registerFile.scala 15:26]
  reg [31:0] _RAND_21;
  reg [31:0] registers_22; // @[registerFile.scala 15:26]
  reg [31:0] _RAND_22;
  reg [31:0] registers_23; // @[registerFile.scala 15:26]
  reg [31:0] _RAND_23;
  reg [31:0] registers_24; // @[registerFile.scala 15:26]
  reg [31:0] _RAND_24;
  reg [31:0] registers_25; // @[registerFile.scala 15:26]
  reg [31:0] _RAND_25;
  reg [31:0] registers_26; // @[registerFile.scala 15:26]
  reg [31:0] _RAND_26;
  reg [31:0] registers_27; // @[registerFile.scala 15:26]
  reg [31:0] _RAND_27;
  reg [31:0] registers_28; // @[registerFile.scala 15:26]
  reg [31:0] _RAND_28;
  reg [31:0] registers_29; // @[registerFile.scala 15:26]
  reg [31:0] _RAND_29;
  reg [31:0] registers_30; // @[registerFile.scala 15:26]
  reg [31:0] _RAND_30;
  reg [31:0] registers_31; // @[registerFile.scala 15:26]
  reg [31:0] _RAND_31;
  wire [31:0] _GEN_1; // @[registerFile.scala 17:10]
  wire [31:0] _GEN_2; // @[registerFile.scala 17:10]
  wire [31:0] _GEN_3; // @[registerFile.scala 17:10]
  wire [31:0] _GEN_4; // @[registerFile.scala 17:10]
  wire [31:0] _GEN_5; // @[registerFile.scala 17:10]
  wire [31:0] _GEN_6; // @[registerFile.scala 17:10]
  wire [31:0] _GEN_7; // @[registerFile.scala 17:10]
  wire [31:0] _GEN_8; // @[registerFile.scala 17:10]
  wire [31:0] _GEN_9; // @[registerFile.scala 17:10]
  wire [31:0] _GEN_10; // @[registerFile.scala 17:10]
  wire [31:0] _GEN_11; // @[registerFile.scala 17:10]
  wire [31:0] _GEN_12; // @[registerFile.scala 17:10]
  wire [31:0] _GEN_13; // @[registerFile.scala 17:10]
  wire [31:0] _GEN_14; // @[registerFile.scala 17:10]
  wire [31:0] _GEN_15; // @[registerFile.scala 17:10]
  wire [31:0] _GEN_16; // @[registerFile.scala 17:10]
  wire [31:0] _GEN_17; // @[registerFile.scala 17:10]
  wire [31:0] _GEN_18; // @[registerFile.scala 17:10]
  wire [31:0] _GEN_19; // @[registerFile.scala 17:10]
  wire [31:0] _GEN_20; // @[registerFile.scala 17:10]
  wire [31:0] _GEN_21; // @[registerFile.scala 17:10]
  wire [31:0] _GEN_22; // @[registerFile.scala 17:10]
  wire [31:0] _GEN_23; // @[registerFile.scala 17:10]
  wire [31:0] _GEN_24; // @[registerFile.scala 17:10]
  wire [31:0] _GEN_25; // @[registerFile.scala 17:10]
  wire [31:0] _GEN_26; // @[registerFile.scala 17:10]
  wire [31:0] _GEN_27; // @[registerFile.scala 17:10]
  wire [31:0] _GEN_28; // @[registerFile.scala 17:10]
  wire [31:0] _GEN_29; // @[registerFile.scala 17:10]
  wire [31:0] _GEN_30; // @[registerFile.scala 17:10]
  wire [31:0] _GEN_33; // @[registerFile.scala 18:10]
  wire [31:0] _GEN_34; // @[registerFile.scala 18:10]
  wire [31:0] _GEN_35; // @[registerFile.scala 18:10]
  wire [31:0] _GEN_36; // @[registerFile.scala 18:10]
  wire [31:0] _GEN_37; // @[registerFile.scala 18:10]
  wire [31:0] _GEN_38; // @[registerFile.scala 18:10]
  wire [31:0] _GEN_39; // @[registerFile.scala 18:10]
  wire [31:0] _GEN_40; // @[registerFile.scala 18:10]
  wire [31:0] _GEN_41; // @[registerFile.scala 18:10]
  wire [31:0] _GEN_42; // @[registerFile.scala 18:10]
  wire [31:0] _GEN_43; // @[registerFile.scala 18:10]
  wire [31:0] _GEN_44; // @[registerFile.scala 18:10]
  wire [31:0] _GEN_45; // @[registerFile.scala 18:10]
  wire [31:0] _GEN_46; // @[registerFile.scala 18:10]
  wire [31:0] _GEN_47; // @[registerFile.scala 18:10]
  wire [31:0] _GEN_48; // @[registerFile.scala 18:10]
  wire [31:0] _GEN_49; // @[registerFile.scala 18:10]
  wire [31:0] _GEN_50; // @[registerFile.scala 18:10]
  wire [31:0] _GEN_51; // @[registerFile.scala 18:10]
  wire [31:0] _GEN_52; // @[registerFile.scala 18:10]
  wire [31:0] _GEN_53; // @[registerFile.scala 18:10]
  wire [31:0] _GEN_54; // @[registerFile.scala 18:10]
  wire [31:0] _GEN_55; // @[registerFile.scala 18:10]
  wire [31:0] _GEN_56; // @[registerFile.scala 18:10]
  wire [31:0] _GEN_57; // @[registerFile.scala 18:10]
  wire [31:0] _GEN_58; // @[registerFile.scala 18:10]
  wire [31:0] _GEN_59; // @[registerFile.scala 18:10]
  wire [31:0] _GEN_60; // @[registerFile.scala 18:10]
  wire [31:0] _GEN_61; // @[registerFile.scala 18:10]
  wire [31:0] _GEN_62; // @[registerFile.scala 18:10]
  wire [31:0] _GEN_64; // @[registerFile.scala 20:26]
  wire [31:0] _GEN_65; // @[registerFile.scala 20:26]
  wire [31:0] _GEN_66; // @[registerFile.scala 20:26]
  wire [31:0] _GEN_67; // @[registerFile.scala 20:26]
  wire [31:0] _GEN_68; // @[registerFile.scala 20:26]
  wire [31:0] _GEN_69; // @[registerFile.scala 20:26]
  wire [31:0] _GEN_70; // @[registerFile.scala 20:26]
  wire [31:0] _GEN_71; // @[registerFile.scala 20:26]
  wire [31:0] _GEN_72; // @[registerFile.scala 20:26]
  wire [31:0] _GEN_73; // @[registerFile.scala 20:26]
  wire [31:0] _GEN_74; // @[registerFile.scala 20:26]
  wire [31:0] _GEN_75; // @[registerFile.scala 20:26]
  wire [31:0] _GEN_76; // @[registerFile.scala 20:26]
  wire [31:0] _GEN_77; // @[registerFile.scala 20:26]
  wire [31:0] _GEN_78; // @[registerFile.scala 20:26]
  wire [31:0] _GEN_79; // @[registerFile.scala 20:26]
  wire [31:0] _GEN_80; // @[registerFile.scala 20:26]
  wire [31:0] _GEN_81; // @[registerFile.scala 20:26]
  wire [31:0] _GEN_82; // @[registerFile.scala 20:26]
  wire [31:0] _GEN_83; // @[registerFile.scala 20:26]
  wire [31:0] _GEN_84; // @[registerFile.scala 20:26]
  wire [31:0] _GEN_85; // @[registerFile.scala 20:26]
  wire [31:0] _GEN_86; // @[registerFile.scala 20:26]
  wire [31:0] _GEN_87; // @[registerFile.scala 20:26]
  wire [31:0] _GEN_88; // @[registerFile.scala 20:26]
  wire [31:0] _GEN_89; // @[registerFile.scala 20:26]
  wire [31:0] _GEN_90; // @[registerFile.scala 20:26]
  wire [31:0] _GEN_91; // @[registerFile.scala 20:26]
  wire [31:0] _GEN_92; // @[registerFile.scala 20:26]
  wire [31:0] _GEN_93; // @[registerFile.scala 20:26]
  wire [31:0] _GEN_94; // @[registerFile.scala 20:26]
  wire [31:0] _GEN_95; // @[registerFile.scala 20:26]
  wire [31:0] _GEN_96; // @[registerFile.scala 19:28]
  wire [31:0] _GEN_97; // @[registerFile.scala 19:28]
  wire [31:0] _GEN_98; // @[registerFile.scala 19:28]
  wire [31:0] _GEN_99; // @[registerFile.scala 19:28]
  wire [31:0] _GEN_100; // @[registerFile.scala 19:28]
  wire [31:0] _GEN_101; // @[registerFile.scala 19:28]
  wire [31:0] _GEN_102; // @[registerFile.scala 19:28]
  wire [31:0] _GEN_103; // @[registerFile.scala 19:28]
  wire [31:0] _GEN_104; // @[registerFile.scala 19:28]
  wire [31:0] _GEN_105; // @[registerFile.scala 19:28]
  wire [31:0] _GEN_106; // @[registerFile.scala 19:28]
  wire [31:0] _GEN_107; // @[registerFile.scala 19:28]
  wire [31:0] _GEN_108; // @[registerFile.scala 19:28]
  wire [31:0] _GEN_109; // @[registerFile.scala 19:28]
  wire [31:0] _GEN_110; // @[registerFile.scala 19:28]
  wire [31:0] _GEN_111; // @[registerFile.scala 19:28]
  wire [31:0] _GEN_112; // @[registerFile.scala 19:28]
  wire [31:0] _GEN_113; // @[registerFile.scala 19:28]
  wire [31:0] _GEN_114; // @[registerFile.scala 19:28]
  wire [31:0] _GEN_115; // @[registerFile.scala 19:28]
  wire [31:0] _GEN_116; // @[registerFile.scala 19:28]
  wire [31:0] _GEN_117; // @[registerFile.scala 19:28]
  wire [31:0] _GEN_118; // @[registerFile.scala 19:28]
  wire [31:0] _GEN_119; // @[registerFile.scala 19:28]
  wire [31:0] _GEN_120; // @[registerFile.scala 19:28]
  wire [31:0] _GEN_121; // @[registerFile.scala 19:28]
  wire [31:0] _GEN_122; // @[registerFile.scala 19:28]
  wire [31:0] _GEN_123; // @[registerFile.scala 19:28]
  wire [31:0] _GEN_124; // @[registerFile.scala 19:28]
  wire [31:0] _GEN_125; // @[registerFile.scala 19:28]
  wire [31:0] _GEN_126; // @[registerFile.scala 19:28]
  wire [31:0] _GEN_127; // @[registerFile.scala 19:28]
  assign _GEN_1 = 5'h1 == io_rs1_sel ? $signed(registers_1) : $signed(registers_0); // @[registerFile.scala 17:10]
  assign _GEN_2 = 5'h2 == io_rs1_sel ? $signed(registers_2) : $signed(_GEN_1); // @[registerFile.scala 17:10]
  assign _GEN_3 = 5'h3 == io_rs1_sel ? $signed(registers_3) : $signed(_GEN_2); // @[registerFile.scala 17:10]
  assign _GEN_4 = 5'h4 == io_rs1_sel ? $signed(registers_4) : $signed(_GEN_3); // @[registerFile.scala 17:10]
  assign _GEN_5 = 5'h5 == io_rs1_sel ? $signed(registers_5) : $signed(_GEN_4); // @[registerFile.scala 17:10]
  assign _GEN_6 = 5'h6 == io_rs1_sel ? $signed(registers_6) : $signed(_GEN_5); // @[registerFile.scala 17:10]
  assign _GEN_7 = 5'h7 == io_rs1_sel ? $signed(registers_7) : $signed(_GEN_6); // @[registerFile.scala 17:10]
  assign _GEN_8 = 5'h8 == io_rs1_sel ? $signed(registers_8) : $signed(_GEN_7); // @[registerFile.scala 17:10]
  assign _GEN_9 = 5'h9 == io_rs1_sel ? $signed(registers_9) : $signed(_GEN_8); // @[registerFile.scala 17:10]
  assign _GEN_10 = 5'ha == io_rs1_sel ? $signed(registers_10) : $signed(_GEN_9); // @[registerFile.scala 17:10]
  assign _GEN_11 = 5'hb == io_rs1_sel ? $signed(registers_11) : $signed(_GEN_10); // @[registerFile.scala 17:10]
  assign _GEN_12 = 5'hc == io_rs1_sel ? $signed(registers_12) : $signed(_GEN_11); // @[registerFile.scala 17:10]
  assign _GEN_13 = 5'hd == io_rs1_sel ? $signed(registers_13) : $signed(_GEN_12); // @[registerFile.scala 17:10]
  assign _GEN_14 = 5'he == io_rs1_sel ? $signed(registers_14) : $signed(_GEN_13); // @[registerFile.scala 17:10]
  assign _GEN_15 = 5'hf == io_rs1_sel ? $signed(registers_15) : $signed(_GEN_14); // @[registerFile.scala 17:10]
  assign _GEN_16 = 5'h10 == io_rs1_sel ? $signed(registers_16) : $signed(_GEN_15); // @[registerFile.scala 17:10]
  assign _GEN_17 = 5'h11 == io_rs1_sel ? $signed(registers_17) : $signed(_GEN_16); // @[registerFile.scala 17:10]
  assign _GEN_18 = 5'h12 == io_rs1_sel ? $signed(registers_18) : $signed(_GEN_17); // @[registerFile.scala 17:10]
  assign _GEN_19 = 5'h13 == io_rs1_sel ? $signed(registers_19) : $signed(_GEN_18); // @[registerFile.scala 17:10]
  assign _GEN_20 = 5'h14 == io_rs1_sel ? $signed(registers_20) : $signed(_GEN_19); // @[registerFile.scala 17:10]
  assign _GEN_21 = 5'h15 == io_rs1_sel ? $signed(registers_21) : $signed(_GEN_20); // @[registerFile.scala 17:10]
  assign _GEN_22 = 5'h16 == io_rs1_sel ? $signed(registers_22) : $signed(_GEN_21); // @[registerFile.scala 17:10]
  assign _GEN_23 = 5'h17 == io_rs1_sel ? $signed(registers_23) : $signed(_GEN_22); // @[registerFile.scala 17:10]
  assign _GEN_24 = 5'h18 == io_rs1_sel ? $signed(registers_24) : $signed(_GEN_23); // @[registerFile.scala 17:10]
  assign _GEN_25 = 5'h19 == io_rs1_sel ? $signed(registers_25) : $signed(_GEN_24); // @[registerFile.scala 17:10]
  assign _GEN_26 = 5'h1a == io_rs1_sel ? $signed(registers_26) : $signed(_GEN_25); // @[registerFile.scala 17:10]
  assign _GEN_27 = 5'h1b == io_rs1_sel ? $signed(registers_27) : $signed(_GEN_26); // @[registerFile.scala 17:10]
  assign _GEN_28 = 5'h1c == io_rs1_sel ? $signed(registers_28) : $signed(_GEN_27); // @[registerFile.scala 17:10]
  assign _GEN_29 = 5'h1d == io_rs1_sel ? $signed(registers_29) : $signed(_GEN_28); // @[registerFile.scala 17:10]
  assign _GEN_30 = 5'h1e == io_rs1_sel ? $signed(registers_30) : $signed(_GEN_29); // @[registerFile.scala 17:10]
  assign _GEN_33 = 5'h1 == io_rs2_sel ? $signed(registers_1) : $signed(registers_0); // @[registerFile.scala 18:10]
  assign _GEN_34 = 5'h2 == io_rs2_sel ? $signed(registers_2) : $signed(_GEN_33); // @[registerFile.scala 18:10]
  assign _GEN_35 = 5'h3 == io_rs2_sel ? $signed(registers_3) : $signed(_GEN_34); // @[registerFile.scala 18:10]
  assign _GEN_36 = 5'h4 == io_rs2_sel ? $signed(registers_4) : $signed(_GEN_35); // @[registerFile.scala 18:10]
  assign _GEN_37 = 5'h5 == io_rs2_sel ? $signed(registers_5) : $signed(_GEN_36); // @[registerFile.scala 18:10]
  assign _GEN_38 = 5'h6 == io_rs2_sel ? $signed(registers_6) : $signed(_GEN_37); // @[registerFile.scala 18:10]
  assign _GEN_39 = 5'h7 == io_rs2_sel ? $signed(registers_7) : $signed(_GEN_38); // @[registerFile.scala 18:10]
  assign _GEN_40 = 5'h8 == io_rs2_sel ? $signed(registers_8) : $signed(_GEN_39); // @[registerFile.scala 18:10]
  assign _GEN_41 = 5'h9 == io_rs2_sel ? $signed(registers_9) : $signed(_GEN_40); // @[registerFile.scala 18:10]
  assign _GEN_42 = 5'ha == io_rs2_sel ? $signed(registers_10) : $signed(_GEN_41); // @[registerFile.scala 18:10]
  assign _GEN_43 = 5'hb == io_rs2_sel ? $signed(registers_11) : $signed(_GEN_42); // @[registerFile.scala 18:10]
  assign _GEN_44 = 5'hc == io_rs2_sel ? $signed(registers_12) : $signed(_GEN_43); // @[registerFile.scala 18:10]
  assign _GEN_45 = 5'hd == io_rs2_sel ? $signed(registers_13) : $signed(_GEN_44); // @[registerFile.scala 18:10]
  assign _GEN_46 = 5'he == io_rs2_sel ? $signed(registers_14) : $signed(_GEN_45); // @[registerFile.scala 18:10]
  assign _GEN_47 = 5'hf == io_rs2_sel ? $signed(registers_15) : $signed(_GEN_46); // @[registerFile.scala 18:10]
  assign _GEN_48 = 5'h10 == io_rs2_sel ? $signed(registers_16) : $signed(_GEN_47); // @[registerFile.scala 18:10]
  assign _GEN_49 = 5'h11 == io_rs2_sel ? $signed(registers_17) : $signed(_GEN_48); // @[registerFile.scala 18:10]
  assign _GEN_50 = 5'h12 == io_rs2_sel ? $signed(registers_18) : $signed(_GEN_49); // @[registerFile.scala 18:10]
  assign _GEN_51 = 5'h13 == io_rs2_sel ? $signed(registers_19) : $signed(_GEN_50); // @[registerFile.scala 18:10]
  assign _GEN_52 = 5'h14 == io_rs2_sel ? $signed(registers_20) : $signed(_GEN_51); // @[registerFile.scala 18:10]
  assign _GEN_53 = 5'h15 == io_rs2_sel ? $signed(registers_21) : $signed(_GEN_52); // @[registerFile.scala 18:10]
  assign _GEN_54 = 5'h16 == io_rs2_sel ? $signed(registers_22) : $signed(_GEN_53); // @[registerFile.scala 18:10]
  assign _GEN_55 = 5'h17 == io_rs2_sel ? $signed(registers_23) : $signed(_GEN_54); // @[registerFile.scala 18:10]
  assign _GEN_56 = 5'h18 == io_rs2_sel ? $signed(registers_24) : $signed(_GEN_55); // @[registerFile.scala 18:10]
  assign _GEN_57 = 5'h19 == io_rs2_sel ? $signed(registers_25) : $signed(_GEN_56); // @[registerFile.scala 18:10]
  assign _GEN_58 = 5'h1a == io_rs2_sel ? $signed(registers_26) : $signed(_GEN_57); // @[registerFile.scala 18:10]
  assign _GEN_59 = 5'h1b == io_rs2_sel ? $signed(registers_27) : $signed(_GEN_58); // @[registerFile.scala 18:10]
  assign _GEN_60 = 5'h1c == io_rs2_sel ? $signed(registers_28) : $signed(_GEN_59); // @[registerFile.scala 18:10]
  assign _GEN_61 = 5'h1d == io_rs2_sel ? $signed(registers_29) : $signed(_GEN_60); // @[registerFile.scala 18:10]
  assign _GEN_62 = 5'h1e == io_rs2_sel ? $signed(registers_30) : $signed(_GEN_61); // @[registerFile.scala 18:10]
  assign _GEN_64 = 5'h0 == io_rd_sel ? $signed(io_writeData) : $signed(32'sh0); // @[registerFile.scala 20:26]
  assign _GEN_65 = 5'h1 == io_rd_sel ? $signed(io_writeData) : $signed(registers_1); // @[registerFile.scala 20:26]
  assign _GEN_66 = 5'h2 == io_rd_sel ? $signed(io_writeData) : $signed(registers_2); // @[registerFile.scala 20:26]
  assign _GEN_67 = 5'h3 == io_rd_sel ? $signed(io_writeData) : $signed(registers_3); // @[registerFile.scala 20:26]
  assign _GEN_68 = 5'h4 == io_rd_sel ? $signed(io_writeData) : $signed(registers_4); // @[registerFile.scala 20:26]
  assign _GEN_69 = 5'h5 == io_rd_sel ? $signed(io_writeData) : $signed(registers_5); // @[registerFile.scala 20:26]
  assign _GEN_70 = 5'h6 == io_rd_sel ? $signed(io_writeData) : $signed(registers_6); // @[registerFile.scala 20:26]
  assign _GEN_71 = 5'h7 == io_rd_sel ? $signed(io_writeData) : $signed(registers_7); // @[registerFile.scala 20:26]
  assign _GEN_72 = 5'h8 == io_rd_sel ? $signed(io_writeData) : $signed(registers_8); // @[registerFile.scala 20:26]
  assign _GEN_73 = 5'h9 == io_rd_sel ? $signed(io_writeData) : $signed(registers_9); // @[registerFile.scala 20:26]
  assign _GEN_74 = 5'ha == io_rd_sel ? $signed(io_writeData) : $signed(registers_10); // @[registerFile.scala 20:26]
  assign _GEN_75 = 5'hb == io_rd_sel ? $signed(io_writeData) : $signed(registers_11); // @[registerFile.scala 20:26]
  assign _GEN_76 = 5'hc == io_rd_sel ? $signed(io_writeData) : $signed(registers_12); // @[registerFile.scala 20:26]
  assign _GEN_77 = 5'hd == io_rd_sel ? $signed(io_writeData) : $signed(registers_13); // @[registerFile.scala 20:26]
  assign _GEN_78 = 5'he == io_rd_sel ? $signed(io_writeData) : $signed(registers_14); // @[registerFile.scala 20:26]
  assign _GEN_79 = 5'hf == io_rd_sel ? $signed(io_writeData) : $signed(registers_15); // @[registerFile.scala 20:26]
  assign _GEN_80 = 5'h10 == io_rd_sel ? $signed(io_writeData) : $signed(registers_16); // @[registerFile.scala 20:26]
  assign _GEN_81 = 5'h11 == io_rd_sel ? $signed(io_writeData) : $signed(registers_17); // @[registerFile.scala 20:26]
  assign _GEN_82 = 5'h12 == io_rd_sel ? $signed(io_writeData) : $signed(registers_18); // @[registerFile.scala 20:26]
  assign _GEN_83 = 5'h13 == io_rd_sel ? $signed(io_writeData) : $signed(registers_19); // @[registerFile.scala 20:26]
  assign _GEN_84 = 5'h14 == io_rd_sel ? $signed(io_writeData) : $signed(registers_20); // @[registerFile.scala 20:26]
  assign _GEN_85 = 5'h15 == io_rd_sel ? $signed(io_writeData) : $signed(registers_21); // @[registerFile.scala 20:26]
  assign _GEN_86 = 5'h16 == io_rd_sel ? $signed(io_writeData) : $signed(registers_22); // @[registerFile.scala 20:26]
  assign _GEN_87 = 5'h17 == io_rd_sel ? $signed(io_writeData) : $signed(registers_23); // @[registerFile.scala 20:26]
  assign _GEN_88 = 5'h18 == io_rd_sel ? $signed(io_writeData) : $signed(registers_24); // @[registerFile.scala 20:26]
  assign _GEN_89 = 5'h19 == io_rd_sel ? $signed(io_writeData) : $signed(registers_25); // @[registerFile.scala 20:26]
  assign _GEN_90 = 5'h1a == io_rd_sel ? $signed(io_writeData) : $signed(registers_26); // @[registerFile.scala 20:26]
  assign _GEN_91 = 5'h1b == io_rd_sel ? $signed(io_writeData) : $signed(registers_27); // @[registerFile.scala 20:26]
  assign _GEN_92 = 5'h1c == io_rd_sel ? $signed(io_writeData) : $signed(registers_28); // @[registerFile.scala 20:26]
  assign _GEN_93 = 5'h1d == io_rd_sel ? $signed(io_writeData) : $signed(registers_29); // @[registerFile.scala 20:26]
  assign _GEN_94 = 5'h1e == io_rd_sel ? $signed(io_writeData) : $signed(registers_30); // @[registerFile.scala 20:26]
  assign _GEN_95 = 5'h1f == io_rd_sel ? $signed(io_writeData) : $signed(registers_31); // @[registerFile.scala 20:26]
  assign _GEN_96 = io_regWrite ? $signed(_GEN_64) : $signed(32'sh0); // @[registerFile.scala 19:28]
  assign _GEN_97 = io_regWrite ? $signed(_GEN_65) : $signed(registers_1); // @[registerFile.scala 19:28]
  assign _GEN_98 = io_regWrite ? $signed(_GEN_66) : $signed(registers_2); // @[registerFile.scala 19:28]
  assign _GEN_99 = io_regWrite ? $signed(_GEN_67) : $signed(registers_3); // @[registerFile.scala 19:28]
  assign _GEN_100 = io_regWrite ? $signed(_GEN_68) : $signed(registers_4); // @[registerFile.scala 19:28]
  assign _GEN_101 = io_regWrite ? $signed(_GEN_69) : $signed(registers_5); // @[registerFile.scala 19:28]
  assign _GEN_102 = io_regWrite ? $signed(_GEN_70) : $signed(registers_6); // @[registerFile.scala 19:28]
  assign _GEN_103 = io_regWrite ? $signed(_GEN_71) : $signed(registers_7); // @[registerFile.scala 19:28]
  assign _GEN_104 = io_regWrite ? $signed(_GEN_72) : $signed(registers_8); // @[registerFile.scala 19:28]
  assign _GEN_105 = io_regWrite ? $signed(_GEN_73) : $signed(registers_9); // @[registerFile.scala 19:28]
  assign _GEN_106 = io_regWrite ? $signed(_GEN_74) : $signed(registers_10); // @[registerFile.scala 19:28]
  assign _GEN_107 = io_regWrite ? $signed(_GEN_75) : $signed(registers_11); // @[registerFile.scala 19:28]
  assign _GEN_108 = io_regWrite ? $signed(_GEN_76) : $signed(registers_12); // @[registerFile.scala 19:28]
  assign _GEN_109 = io_regWrite ? $signed(_GEN_77) : $signed(registers_13); // @[registerFile.scala 19:28]
  assign _GEN_110 = io_regWrite ? $signed(_GEN_78) : $signed(registers_14); // @[registerFile.scala 19:28]
  assign _GEN_111 = io_regWrite ? $signed(_GEN_79) : $signed(registers_15); // @[registerFile.scala 19:28]
  assign _GEN_112 = io_regWrite ? $signed(_GEN_80) : $signed(registers_16); // @[registerFile.scala 19:28]
  assign _GEN_113 = io_regWrite ? $signed(_GEN_81) : $signed(registers_17); // @[registerFile.scala 19:28]
  assign _GEN_114 = io_regWrite ? $signed(_GEN_82) : $signed(registers_18); // @[registerFile.scala 19:28]
  assign _GEN_115 = io_regWrite ? $signed(_GEN_83) : $signed(registers_19); // @[registerFile.scala 19:28]
  assign _GEN_116 = io_regWrite ? $signed(_GEN_84) : $signed(registers_20); // @[registerFile.scala 19:28]
  assign _GEN_117 = io_regWrite ? $signed(_GEN_85) : $signed(registers_21); // @[registerFile.scala 19:28]
  assign _GEN_118 = io_regWrite ? $signed(_GEN_86) : $signed(registers_22); // @[registerFile.scala 19:28]
  assign _GEN_119 = io_regWrite ? $signed(_GEN_87) : $signed(registers_23); // @[registerFile.scala 19:28]
  assign _GEN_120 = io_regWrite ? $signed(_GEN_88) : $signed(registers_24); // @[registerFile.scala 19:28]
  assign _GEN_121 = io_regWrite ? $signed(_GEN_89) : $signed(registers_25); // @[registerFile.scala 19:28]
  assign _GEN_122 = io_regWrite ? $signed(_GEN_90) : $signed(registers_26); // @[registerFile.scala 19:28]
  assign _GEN_123 = io_regWrite ? $signed(_GEN_91) : $signed(registers_27); // @[registerFile.scala 19:28]
  assign _GEN_124 = io_regWrite ? $signed(_GEN_92) : $signed(registers_28); // @[registerFile.scala 19:28]
  assign _GEN_125 = io_regWrite ? $signed(_GEN_93) : $signed(registers_29); // @[registerFile.scala 19:28]
  assign _GEN_126 = io_regWrite ? $signed(_GEN_94) : $signed(registers_30); // @[registerFile.scala 19:28]
  assign _GEN_127 = io_regWrite ? $signed(_GEN_95) : $signed(registers_31); // @[registerFile.scala 19:28]
  assign io_rs1 = 5'h1f == io_rs1_sel ? $signed(registers_31) : $signed(_GEN_30); // @[registerFile.scala 17:10]
  assign io_rs2 = 5'h1f == io_rs2_sel ? $signed(registers_31) : $signed(_GEN_62); // @[registerFile.scala 18:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  registers_0 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  registers_1 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  registers_2 = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  registers_3 = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  registers_4 = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  registers_5 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  registers_6 = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  registers_7 = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  registers_8 = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  registers_9 = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  registers_10 = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  registers_11 = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  registers_12 = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  registers_13 = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  registers_14 = _RAND_14[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  registers_15 = _RAND_15[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  registers_16 = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  registers_17 = _RAND_17[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  registers_18 = _RAND_18[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  registers_19 = _RAND_19[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  registers_20 = _RAND_20[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  registers_21 = _RAND_21[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  registers_22 = _RAND_22[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  registers_23 = _RAND_23[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  registers_24 = _RAND_24[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  registers_25 = _RAND_25[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  registers_26 = _RAND_26[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  registers_27 = _RAND_27[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  registers_28 = _RAND_28[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  registers_29 = _RAND_29[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  registers_30 = _RAND_30[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  registers_31 = _RAND_31[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      registers_0 <= 32'sh0;
    end else begin
      if (io_regWrite) begin
        if (5'h0 == io_rd_sel) begin
          registers_0 <= io_writeData;
        end else begin
          registers_0 <= 32'sh0;
        end
      end else begin
        registers_0 <= 32'sh0;
      end
    end
    if (reset) begin
      registers_1 <= 32'sh0;
    end else begin
      if (io_regWrite) begin
        if (5'h1 == io_rd_sel) begin
          registers_1 <= io_writeData;
        end
      end
    end
    if (reset) begin
      registers_2 <= 32'sh0;
    end else begin
      if (io_regWrite) begin
        if (5'h2 == io_rd_sel) begin
          registers_2 <= io_writeData;
        end
      end
    end
    if (reset) begin
      registers_3 <= 32'sh0;
    end else begin
      if (io_regWrite) begin
        if (5'h3 == io_rd_sel) begin
          registers_3 <= io_writeData;
        end
      end
    end
    if (reset) begin
      registers_4 <= 32'sh0;
    end else begin
      if (io_regWrite) begin
        if (5'h4 == io_rd_sel) begin
          registers_4 <= io_writeData;
        end
      end
    end
    if (reset) begin
      registers_5 <= 32'sh0;
    end else begin
      if (io_regWrite) begin
        if (5'h5 == io_rd_sel) begin
          registers_5 <= io_writeData;
        end
      end
    end
    if (reset) begin
      registers_6 <= 32'sh0;
    end else begin
      if (io_regWrite) begin
        if (5'h6 == io_rd_sel) begin
          registers_6 <= io_writeData;
        end
      end
    end
    if (reset) begin
      registers_7 <= 32'sh0;
    end else begin
      if (io_regWrite) begin
        if (5'h7 == io_rd_sel) begin
          registers_7 <= io_writeData;
        end
      end
    end
    if (reset) begin
      registers_8 <= 32'sh0;
    end else begin
      if (io_regWrite) begin
        if (5'h8 == io_rd_sel) begin
          registers_8 <= io_writeData;
        end
      end
    end
    if (reset) begin
      registers_9 <= 32'sh0;
    end else begin
      if (io_regWrite) begin
        if (5'h9 == io_rd_sel) begin
          registers_9 <= io_writeData;
        end
      end
    end
    if (reset) begin
      registers_10 <= 32'sh0;
    end else begin
      if (io_regWrite) begin
        if (5'ha == io_rd_sel) begin
          registers_10 <= io_writeData;
        end
      end
    end
    if (reset) begin
      registers_11 <= 32'sh0;
    end else begin
      if (io_regWrite) begin
        if (5'hb == io_rd_sel) begin
          registers_11 <= io_writeData;
        end
      end
    end
    if (reset) begin
      registers_12 <= 32'sh0;
    end else begin
      if (io_regWrite) begin
        if (5'hc == io_rd_sel) begin
          registers_12 <= io_writeData;
        end
      end
    end
    if (reset) begin
      registers_13 <= 32'sh0;
    end else begin
      if (io_regWrite) begin
        if (5'hd == io_rd_sel) begin
          registers_13 <= io_writeData;
        end
      end
    end
    if (reset) begin
      registers_14 <= 32'sh0;
    end else begin
      if (io_regWrite) begin
        if (5'he == io_rd_sel) begin
          registers_14 <= io_writeData;
        end
      end
    end
    if (reset) begin
      registers_15 <= 32'sh0;
    end else begin
      if (io_regWrite) begin
        if (5'hf == io_rd_sel) begin
          registers_15 <= io_writeData;
        end
      end
    end
    if (reset) begin
      registers_16 <= 32'sh0;
    end else begin
      if (io_regWrite) begin
        if (5'h10 == io_rd_sel) begin
          registers_16 <= io_writeData;
        end
      end
    end
    if (reset) begin
      registers_17 <= 32'sh0;
    end else begin
      if (io_regWrite) begin
        if (5'h11 == io_rd_sel) begin
          registers_17 <= io_writeData;
        end
      end
    end
    if (reset) begin
      registers_18 <= 32'sh0;
    end else begin
      if (io_regWrite) begin
        if (5'h12 == io_rd_sel) begin
          registers_18 <= io_writeData;
        end
      end
    end
    if (reset) begin
      registers_19 <= 32'sh0;
    end else begin
      if (io_regWrite) begin
        if (5'h13 == io_rd_sel) begin
          registers_19 <= io_writeData;
        end
      end
    end
    if (reset) begin
      registers_20 <= 32'sh0;
    end else begin
      if (io_regWrite) begin
        if (5'h14 == io_rd_sel) begin
          registers_20 <= io_writeData;
        end
      end
    end
    if (reset) begin
      registers_21 <= 32'sh0;
    end else begin
      if (io_regWrite) begin
        if (5'h15 == io_rd_sel) begin
          registers_21 <= io_writeData;
        end
      end
    end
    if (reset) begin
      registers_22 <= 32'sh0;
    end else begin
      if (io_regWrite) begin
        if (5'h16 == io_rd_sel) begin
          registers_22 <= io_writeData;
        end
      end
    end
    if (reset) begin
      registers_23 <= 32'sh0;
    end else begin
      if (io_regWrite) begin
        if (5'h17 == io_rd_sel) begin
          registers_23 <= io_writeData;
        end
      end
    end
    if (reset) begin
      registers_24 <= 32'sh0;
    end else begin
      if (io_regWrite) begin
        if (5'h18 == io_rd_sel) begin
          registers_24 <= io_writeData;
        end
      end
    end
    if (reset) begin
      registers_25 <= 32'sh0;
    end else begin
      if (io_regWrite) begin
        if (5'h19 == io_rd_sel) begin
          registers_25 <= io_writeData;
        end
      end
    end
    if (reset) begin
      registers_26 <= 32'sh0;
    end else begin
      if (io_regWrite) begin
        if (5'h1a == io_rd_sel) begin
          registers_26 <= io_writeData;
        end
      end
    end
    if (reset) begin
      registers_27 <= 32'sh0;
    end else begin
      if (io_regWrite) begin
        if (5'h1b == io_rd_sel) begin
          registers_27 <= io_writeData;
        end
      end
    end
    if (reset) begin
      registers_28 <= 32'sh0;
    end else begin
      if (io_regWrite) begin
        if (5'h1c == io_rd_sel) begin
          registers_28 <= io_writeData;
        end
      end
    end
    if (reset) begin
      registers_29 <= 32'sh0;
    end else begin
      if (io_regWrite) begin
        if (5'h1d == io_rd_sel) begin
          registers_29 <= io_writeData;
        end
      end
    end
    if (reset) begin
      registers_30 <= 32'sh0;
    end else begin
      if (io_regWrite) begin
        if (5'h1e == io_rd_sel) begin
          registers_30 <= io_writeData;
        end
      end
    end
    if (reset) begin
      registers_31 <= 32'sh0;
    end else begin
      if (io_regWrite) begin
        if (5'h1f == io_rd_sel) begin
          registers_31 <= io_writeData;
        end
      end
    end
  end
endmodule
